module hexdriver (input [3:0] val, output logic [6:0] hex);
    /*
    * if 0000
    * output 7'b0000001
    * elif 0001
    * ...
    * elif 1001
    */
    assign hex = 
        val == 4'b0000 ? 7'b1000000 : // 0
        val == 4'b0001 ? 7'b1111001 : // 1
        val == 4'b0010 ? 7'b0100100 : // 2
        val == 4'b0011 ? 7'b0110000 : // 3
        val == 4'b0100 ? 7'b0011001 : // 4
        val == 4'b0101 ? 7'b0010010 : // 5
        val == 4'b0110 ? 7'b0000010 : // 6
        val == 4'b0111 ? 7'b1111000 : // 7
        val == 4'b1000 ? 7'b0000000 : // 8
        val == 4'b1001 ? 7'b0010000 : // 9
        val == 4'b1010 ? 7'b0001000 : // 10 (A)
        val == 4'b1011 ? 7'b0000011 : // 11 (b)
        val == 4'b1100 ? 7'b1000110 : // 12 (C)
        val == 4'b1101 ? 7'b0100001 : // 13 (d)
        val == 4'b1110 ? 7'b0000110 : // 14 (E)
        val == 4'b1111 ? 7'b0001110 : // 15 (F)

           7'b0111111;	     // default (error case)
endmodule
